----------------------------------------------------------------------------------
-- Company: N/A
-- Engineer: Kyle Gapinski
-- 
-- Create Date:    12:48:11 02/01/2016 
-- Design Name: IDR Virtualization
-- Module Name:    Top_Module - Behavioral 
-- Project Name: Capstone Project
-- Target Devices: Unknown 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Top_Module is
end Top_Module;

architecture Behavioral of Top_Module is

begin
--This is place holder for future project.

end Behavioral;

